�� 
 / /   C o d e   y o u r   d e s i g n   h e r e  
 ` t i m e s c a l e   1 n s   /   1 p s  
  
 m o d u l e   R I S C _ S P M   ( c l k ,   r s t ,   a l u _ o u t _ t e m p e r a t u r e ,   a l u _ o u t _ b a t t e r y ,   a l u _ o u t _ G A S ,   a l u _ o u t _ T r a n s m i s s i o n , a l u _ o u t _ P r e s s u r e ,   a l u _ o u t _ O I L ) ;  
     p a r a m e t e r   w o r d _ s i z e   =   9 ;  
     p a r a m e t e r   S e l 1 _ s i z e   =   3 ;  
     p a r a m e t e r   S e l 2 _ s i z e   =   2 ;  
     w i r e   [ S e l 1 _ s i z e - 1 :   0 ]   S e l _ B u s _ 1 _ M u x ;  
     w i r e   [ S e l 2 _ s i z e - 1 :   0 ]   S e l _ B u s _ 2 _ M u x ;  
  
     i n p u t   c l k ,   r s t ;  
  
     / /   D a t a   N e t s  
     w i r e   z e r o ;  
     w i r e   [ w o r d _ s i z e - 1 :   0 ]   i n s t r u c t i o n ,   a d d r e s s ,   B u s _ 1 ,   m e m _ w o r d ;  
        
     / /   C o n t r o l   N e t s  
     w i r e   L o a d _ R 0 ,   L o a d _ R 1 ,   L o a d _ R 2 ,   L o a d _ R 3 ,   L o a d _ P C ,   I n c _ P C ,   L o a d _ I R ;        
     w i r e   L o a d _ A d d _ R ,   L o a d _ R e g _ Y ,   L o a d _ R e g _ Z ;  
     w i r e   w r i t e ;  
   o u t p u t   a l u _ o u t _ t e m p e r a t u r e ,   a l u _ o u t _ b a t t e r y ,   a l u _ o u t _ G A S ,   a l u _ o u t _ T r a n s m i s s i o n , a l u _ o u t _ P r e s s u r e ,   a l u _ o u t _ O I L ;  
    
     P r o c e s s i n g _ U n i t   M 0 _ P r o c e s s o r   ( i n s t r u c t i o n ,   z e r o ,   a d d r e s s ,   B u s _ 1 ,   m e m _ w o r d ,   L o a d _ R 0 ,   L o a d _ R 1 ,  
         L o a d _ R 2 ,   L o a d _ R 3 ,   L o a d _ P C ,   I n c _ P C ,   S e l _ B u s _ 1 _ M u x ,   L o a d _ I R ,   L o a d _ A d d _ R ,   L o a d _ R e g _ Y ,  
         L o a d _ R e g _ Z ,     S e l _ B u s _ 2 _ M u x ,   c l k ,   r s t ,   a l u _ o u t _ t e m p e r a t u r e ,   a l u _ o u t _ b a t t e r y ,   a l u _ o u t _ G A S ,   a l u _ o u t _ T r a n s m i s s i o n , a l u _ o u t _ P r e s s u r e ,   a l u _ o u t _ O I L ) ;  
  
     C o n t r o l _ U n i t   M 1 _ C o n t r o l l e r   ( L o a d _ R 0 ,   L o a d _ R 1 ,   L o a d _ R 2 ,   L o a d _ R 3 ,   L o a d _ P C ,   I n c _ P C ,    
         S e l _ B u s _ 1 _ M u x ,   S e l _ B u s _ 2 _ M u x   ,   L o a d _ I R ,   L o a d _ A d d _ R ,   L o a d _ R e g _ Y ,   L o a d _ R e g _ Z ,    
         w r i t e ,   i n s t r u c t i o n ,   z e r o ,   c l k ,   r s t ) ;  
  
     M e m o r y _ U n i t   M 2 _ S R A M   (  
         . d a t a _ o u t ( m e m _ w o r d ) ,    
         . d a t a _ i n ( B u s _ 1 ) ,    
         . a d d r e s s ( a d d r e s s ) ,    
         . c l k ( c l k ) ,  
         . w r i t e ( w r i t e )   ) ;  
 e n d m o d u l e  
  
  
 m o d u l e   P r o c e s s i n g _ U n i t   ( i n s t r u c t i o n ,   Z f l a g ,   a d d r e s s ,   B u s _ 1 ,   m e m _ w o r d ,   L o a d _ R 0 ,   L o a d _ R 1 ,   L o a d _ R 2 ,    
     L o a d _ R 3 ,   L o a d _ P C ,   I n c _ P C ,   S e l _ B u s _ 1 _ M u x ,   L o a d _ I R ,   L o a d _ A d d _ R ,   L o a d _ R e g _ Y ,   L o a d _ R e g _ Z ,    
     S e l _ B u s _ 2 _ M u x ,   c l k ,   r s t , a l u _ o u t _ t e m p e r a t u r e ,   a l u _ o u t _ b a t t e r y ,   a l u _ o u t _ G A S ,   a l u _ o u t _ T r a n s m i s s i o n , a l u _ o u t _ P r e s s u r e ,   a l u _ o u t _ O I L ) ;  
  
     p a r a m e t e r   w o r d _ s i z e   =   9 ;  
     p a r a m e t e r   o p _ s i z e   =   4 ;  
     p a r a m e t e r   S e l 1 _ s i z e   =   3 ;  
     p a r a m e t e r   S e l 2 _ s i z e   =   2 ;  
  
     o u t p u t   [ w o r d _ s i z e - 1 :   0 ]   	 i n s t r u c t i o n ,   a d d r e s s ,   B u s _ 1 ;  
     o u t p u t   Z f l a g ;  
         o u t p u t     a l u _ o u t _ t e m p e r a t u r e ,   a l u _ o u t _ b a t t e r y ,   a l u _ o u t _ G A S ,   a l u _ o u t _ T r a n s m i s s i o n , a l u _ o u t _ P r e s s u r e ,   a l u _ o u t _ O I L ;  
     i n p u t   [ w o r d _ s i z e - 1 :   0 ]     	 m e m _ w o r d ;  
     i n p u t   	 	 	 L o a d _ R 0 ,   L o a d _ R 1 ,   L o a d _ R 2 ,   L o a d _ R 3 ,   L o a d _ P C ,   I n c _ P C ;  
     i n p u t   [ S e l 1 _ s i z e - 1 :   0 ]   	 S e l _ B u s _ 1 _ M u x ;  
     i n p u t   [ S e l 2 _ s i z e - 1 :   0 ]   	 S e l _ B u s _ 2 _ M u x ;  
     i n p u t   	 	 	 L o a d _ I R ,   L o a d _ A d d _ R ,   L o a d _ R e g _ Y ,   L o a d _ R e g _ Z ;  
     i n p u t   	 	 	 c l k ,   r s t ;  
  
     w i r e 	 	 	 L o a d _ R 0 ,   L o a d _ R 1 ,   L o a d _ R 2 ,   L o a d _ R 3 ;  
     w i r e   [ w o r d _ s i z e - 1 :   0 ]   	 B u s _ 2 ;  
     w i r e   [ w o r d _ s i z e - 1 :   0 ]   	 R 0 _ o u t ,   R 1 _ o u t ,   R 2 _ o u t ,   R 3 _ o u t ;  
     w i r e   [ w o r d _ s i z e - 1 :   0 ]   	 P C _ c o u n t ,   Y _ v a l u e ,   a l u _ o u t ;  
     w i r e   	 	 	 a l u _ z e r o _ f l a g ;  
     w i r e   [ o p _ s i z e - 1   :   0 ]   	 o p c o d e   =   i n s t r u c t i o n   [ w o r d _ s i z e - 1 :   w o r d _ s i z e - o p _ s i z e ] ;  
  
     R e g i s t e r _ U n i t   	 	 R 0   	 ( R 0 _ o u t ,   B u s _ 2 ,   L o a d _ R 0 ,   c l k ,   r s t ) ;  
     R e g i s t e r _ U n i t   	 	 R 1   	 ( R 1 _ o u t ,   B u s _ 2 ,   L o a d _ R 1 ,   c l k ,   r s t ) ;  
     R e g i s t e r _ U n i t   	 	 R 2   	 ( R 2 _ o u t ,   B u s _ 2 ,   L o a d _ R 2 ,   c l k ,   r s t ) ;  
     R e g i s t e r _ U n i t   	 	 R 3   	 ( R 3 _ o u t ,   B u s _ 2 ,   L o a d _ R 3 ,   c l k ,   r s t ) ;  
     R e g i s t e r _ U n i t   	 	 R e g _ Y   	 ( Y _ v a l u e ,   B u s _ 2 ,   L o a d _ R e g _ Y ,   c l k ,   r s t ) ;  
     D _ f l o p   	 	 	 R e g _ Z   	 ( Z f l a g ,   a l u _ z e r o _ f l a g ,   L o a d _ R e g _ Z ,   c l k ,   r s t ) ;  
     A d d r e s s _ R e g i s t e r   	 A d d _ R 	 ( a d d r e s s ,   B u s _ 2 ,   L o a d _ A d d _ R ,   c l k ,   r s t ) ;  
     I n s t r u c t i o n _ R e g i s t e r 	 I R 	 ( i n s t r u c t i o n ,   B u s _ 2 ,   L o a d _ I R ,   c l k ,   r s t ) ;  
     P r o g r a m _ C o u n t e r   	 P C 	 ( P C _ c o u n t ,   B u s _ 2 ,   L o a d _ P C ,   I n c _ P C ,   c l k ,   r s t ) ;  
     M u l t i p l e x e r _ 5 c h   	 	 M u x _ 1   	 ( B u s _ 1 ,   R 0 _ o u t ,   R 1 _ o u t ,   R 2 _ o u t ,   R 3 _ o u t ,   P C _ c o u n t ,   S e l _ B u s _ 1 _ M u x ) ;  
     M u l t i p l e x e r _ 3 c h   	 	 M u x _ 2 	 ( B u s _ 2 ,   a l u _ o u t ,   B u s _ 1 ,   m e m _ w o r d ,   S e l _ B u s _ 2 _ M u x ) ;  
     A l u _ R I S C   	 	 A L U 	 ( a l u _ z e r o _ f l a g ,   a l u _ o u t ,   Y _ v a l u e ,   B u s _ 1 ,   o p c o d e , a l u _ o u t _ t e m p e r a t u r e ,   a l u _ o u t _ b a t t e r y ,   a l u _ o u t _ G A S ,   a l u _ o u t _ T r a n s m i s s i o n , a l u _ o u t _ P r e s s u r e ,   a l u _ o u t _ O I L ) ;  
 e n d m o d u l e    
  
 m o d u l e   R e g i s t e r _ U n i t   ( d a t a _ o u t ,   d a t a _ i n ,   l o a d ,   c l k ,   r s t ) ;  
     p a r a m e t e r   	 	 w o r d _ s i z e   =   9 ;  
     o u t p u t   [ w o r d _ s i z e - 1 :   0 ]   	 d a t a _ o u t ;  
     i n p u t   	 [ w o r d _ s i z e - 1 :   0 ]   	 d a t a _ i n ;  
     i n p u t   	 	 	 l o a d ;  
     i n p u t   	 	 	 c l k ,   r s t ;  
     r e g   	 [ w o r d _ s i z e - 1 :   0 ] 	 d a t a _ o u t ;  
  
     a l w a y s   @   ( p o s e d g e   c l k   o r   n e g e d g e   r s t )  
         i f   ( r s t   = =   0 )   d a t a _ o u t   < =   0 ;   e l s e   i f   ( l o a d )   d a t a _ o u t   < =   d a t a _ i n ;  
 e n d m o d u l e  
  
 m o d u l e   D _ f l o p   ( d a t a _ o u t ,   d a t a _ i n ,   l o a d ,   c l k ,   r s t ) ;  
     o u t p u t   	 	 d a t a _ o u t ;  
     i n p u t   	 	 d a t a _ i n ;  
     i n p u t   	 	 l o a d ;  
     i n p u t   	 	 c l k ,   r s t ;  
     r e g   	 	 d a t a _ o u t ;  
  
     a l w a y s   @   ( p o s e d g e   c l k   o r   n e g e d g e   r s t )  
         i f   ( r s t   = =   0 )   d a t a _ o u t   < =   0 ;   e l s e   i f   ( l o a d   = =   1 ) d a t a _ o u t   < =   d a t a _ i n ;  
 e n d m o d u l e  
  
   m o d u l e   A d d r e s s _ R e g i s t e r   ( d a t a _ o u t ,   d a t a _ i n ,   l o a d ,   c l k ,   r s t ) ;  
     p a r a m e t e r   w o r d _ s i z e   =   9 ;  
     o u t p u t   [ w o r d _ s i z e - 1 :   0 ]   	 d a t a _ o u t ;  
     i n p u t   	 [ w o r d _ s i z e - 1 :   0 ]   	 d a t a _ i n ;  
     i n p u t   	 	 	 l o a d ,   c l k ,   r s t ;  
     r e g   	 [ w o r d _ s i z e - 1 :   0 ] 	 d a t a _ o u t ;  
     a l w a y s   @   ( p o s e d g e   c l k   o r   n e g e d g e   r s t )  
         i f   ( r s t   = =   0 )   d a t a _ o u t   < =   0 ;   e l s e   i f   ( l o a d )   d a t a _ o u t   < =   d a t a _ i n ;  
 e n d m o d u l e  
  
 m o d u l e   I n s t r u c t i o n _ R e g i s t e r   ( d a t a _ o u t ,   d a t a _ i n ,   l o a d ,   c l k ,   r s t ) ;  
     p a r a m e t e r   w o r d _ s i z e   =   9 ;  
     o u t p u t   [ w o r d _ s i z e - 1 :   0 ]   	 d a t a _ o u t ;  
     i n p u t   	 [ w o r d _ s i z e - 1 :   0 ]   	 d a t a _ i n ;  
     i n p u t   	 	 	 l o a d ;  
     i n p u t   	 	 	 c l k ,   r s t ;  
     r e g   	 [ w o r d _ s i z e - 1 :   0 ] 	 d a t a _ o u t ;  
     a l w a y s   @   ( p o s e d g e   c l k   o r   n e g e d g e   r s t )  
         i f   ( r s t   = =   0 )   d a t a _ o u t   < =   0 ;   e l s e   i f   ( l o a d )   d a t a _ o u t   < =   d a t a _ i n ;    
 e n d m o d u l e  
  
 m o d u l e   P r o g r a m _ C o u n t e r   ( c o u n t ,   d a t a _ i n ,   L o a d _ P C ,   I n c _ P C ,   c l k ,   r s t ) ;  
     p a r a m e t e r   w o r d _ s i z e   =   9 ;  
     o u t p u t   [ w o r d _ s i z e - 1 :   0 ]   	 c o u n t ;  
     i n p u t   	 [ w o r d _ s i z e - 1 :   0 ]   	 d a t a _ i n ;  
     i n p u t   	 	 	 L o a d _ P C ,   I n c _ P C ;  
     i n p u t   	 	 	 c l k ,   r s t ;  
     r e g   	 [ w o r d _ s i z e - 1 :   0 ] 	 c o u n t ;  
     a l w a y s   @   ( p o s e d g e   c l k   o r   n e g e d g e   r s t )  
         i f   ( r s t   = =   0 )   c o u n t   < =   0 ;   e l s e   i f   ( L o a d _ P C )   c o u n t   < =   d a t a _ i n ;   e l s e   i f     ( I n c _ P C )   c o u n t   < =   c o u n t   + 1 ;  
 e n d m o d u l e  
  
 m o d u l e   M u l t i p l e x e r _ 5 c h   ( m u x _ o u t ,   d a t a _ a ,   d a t a _ b ,   d a t a _ c ,   d a t a _ d ,   d a t a _ e ,   s e l ) ;  
     p a r a m e t e r   w o r d _ s i z e   =   9 ;  
     o u t p u t   [ w o r d _ s i z e - 1 :   0 ]   	 m u x _ o u t ;  
     i n p u t   	 [ w o r d _ s i z e - 1 :   0 ]   	 d a t a _ a ,   d a t a _ b ,   d a t a _ c ,   d a t a _ d ,   d a t a _ e ;  
     i n p u t   	 [ 2 :   0 ]   s e l ;  
    
     a s s i g n     m u x _ o u t   =   ( s e l   = =   0 )   	 ?   d a t a _ a :   ( s e l   = =   1 )    
 ?   d a t a _ b   :   ( s e l   = =   2 )    
 ?   d a t a _ c :   ( s e l   = =   3 )    
 ?   d a t a _ d   :   ( s e l   = =   4 )    
 ?   d a t a _ e   :   ' b x ;  
 e n d m o d u l e  
  
 m o d u l e   M u l t i p l e x e r _ 3 c h   ( m u x _ o u t ,   d a t a _ a ,   d a t a _ b ,   d a t a _ c ,   s e l ) ;  
     p a r a m e t e r   	 w o r d _ s i z e   =   9 ;  
     o u t p u t   	 	 [ w o r d _ s i z e - 1 :   0 ] 	   m u x _ o u t ;  
     i n p u t   	 	 [ w o r d _ s i z e - 1 :   0 ]   	 d a t a _ a ,   d a t a _ b ,   d a t a _ c ;  
     i n p u t   	 	 [ 1 :   0 ]   s e l ;  
  
     a s s i g n     m u x _ o u t   =   ( s e l   = =   0 )   ?   d a t a _ a :   ( s e l   = =   1 )   ?   d a t a _ b   :   ( s e l   = =   2 )   ?   d a t a _ c :   ' b x ;  
 e n d m o d u l e  
    
  
  
 / * A L U   I n s t r u c t i o n 	 	 A c t i o n  
 A D D 	 	 	 A d d s   t h e   d a t a p a t h s   t o   f o r m   d a t a _ 1   +   d a t a _ 2 .  
 S U B 	 	 	 S u b t r a c t s   t h e   d a t a p a t h s   t o   f o r m   d a t a _ 1   -   d a t a _ 2 .  
 A N D 	 	 	 T a k e s   t h e   b i t w i s e - a n d   o f   t h e   d a t a p a t h s ,   d a t a _ 1   &   d a t a _ 2 .  
 N O T 	 	 	 T a k e s   t h e   b i t w i s e   B o o l e a n   c o m p l e m e n t   o f   d a t a _ 1 .  
 * /  
 / /   N o t e :   t h e   c a r r i e s   a r e   i g n o r e d   i n   t h i s   m o d e l .  
    
 m o d u l e   A l u _ R I S C   ( a l u _ z e r o _ f l a g ,   a l u _ o u t ,   d a t a _ 1 ,   d a t a _ 2 ,   s e l , a l u _ o u t _ t e m p e r a t u r e ,   a l u _ o u t _ b a t t e r y ,   a l u _ o u t _ G A S ,   a l u _ o u t _ T r a n s m i s s i o n , a l u _ o u t _ P r e s s u r e ,   a l u _ o u t _ O I L ) ;  
     p a r a m e t e r   w o r d _ s i z e   =   9 ;  
     p a r a m e t e r   o p _ s i z e   =   4 ;  
     / /   O p c o d e s  
     p a r a m e t e r   N O P   =   4 ' b 0 0 0 0 ;  
     p a r a m e t e r   A D D   =   4 ' b 0 0 0 1 ;  
     p a r a m e t e r   S U B   =   4 ' b 0 0 1 0 ;  
     p a r a m e t e r   A N D   =   4 ' b 0 0 1 1 ;  
     p a r a m e t e r   N O T   =   4 ' b 0 1 0 0 ;  
     p a r a m e t e r   R D       =   4 ' b 0 1 0 1 ;  
     p a r a m e t e r   W R   =   4 ' b 0 1 1 0 ;  
     p a r a m e t e r   B R   =   4 ' b 0 1 1 1 ;  
     p a r a m e t e r   B R Z   =   4 ' b 1 0 0 0 ;  
    
     p a r a m e t e r   C M P _ G A S           =   4 ' b 1 0 0 1 ;  
     p a r a m e t e r   C M P _ T r a n s m i s s i o n           =   4 ' b 1 0 1 0 ;  
     p a r a m e t e r   C M P _ P r e s s u r e           =   4 ' b 1 0 1 1 ;  
     p a r a m e t e r   C M P _ O I L           =   4 ' b 1 1 0 0 ;  
     p a r a m e t e r   C M P _ T e m p e r a t u r e           =   4 ' b 1 1 0 1 ;  
     p a r a m e t e r   C M P _ b a t t e r y           =   4 ' b 1 1 1 0 ;  
  
     o u t p u t   a l u _ z e r o _ f l a g ;  
     o u t p u t   [ w o r d _ s i z e - 1 :   0 ]   a l u _ o u t ;  
     o u t p u t   r e g   a l u _ o u t _ t e m p e r a t u r e ,   a l u _ o u t _ b a t t e r y ,   a l u _ o u t _ G A S ,   a l u _ o u t _ T r a n s m i s s i o n , a l u _ o u t _ P r e s s u r e ,   a l u _ o u t _ O I L ;  
     i n p u t       [ w o r d _ s i z e - 1 :   0 ]   d a t a _ 1 ,   d a t a _ 2 ;  
     i n p u t   [ o p _ s i z e - 1 :   0 ]   s e l ;  
     r e g   [ w o r d _ s i z e - 1 :   0 ]   a l u _ o u t ;  
      
     i n i t i a l  
     b e g i n  
     a l u _ o u t _ t e m p e r a t u r e   = 0 ;   a l u _ o u t _ b a t t e r y = 0 ;   a l u _ o u t _ G A S   = 0   ; a l u _ o u t _ T r a n s m i s s i o n   = 0 ;  
     a l u _ o u t _ P r e s s u r e = 0 ;   a l u _ o u t _ O I L = 0 ;  
     a l u _ o u t   =   0 ;    
     e n d  
      
  
     a s s i g n     a l u _ z e r o _ f l a g   =   ~ | a l u _ o u t ;  
     a l w a y s   @   ( s e l   o r   d a t a _ 1   o r   d a t a _ 2 )      
           c a s e     ( s e l )  
             N O P :   a l u _ o u t   =   0 ;  
             A D D :   a l u _ o u t   =   d a t a _ 1   +   d a t a _ 2 ;     / /   R e g _ Y   +   B u s _ 1  
             S U B :   a l u _ o u t   =   d a t a _ 2   -   d a t a _ 1 ;  
             A N D :   a l u _ o u t   =   d a t a _ 1   &   d a t a _ 2 ;  
             N O T :   a l u _ o u t   =   ~   d a t a _ 2 ;   / /   G e t s   d a t a   f r o m   B u s _ 1  
            
            
             C M P _ G A S :     i f ( d a t a _ 2 < = 9 ' h 0 f 0 )   b e g i n   a l u _ o u t _ G A S   < =   0 ;   e n d  
                                 e l s e   b e g i n   a l u _ o u t _ G A S   < =   1 ;   e n d  
             C M P _ T r a n s m i s s i o n :     i f ( d a t a _ 2 < = 9 ' h 0 f 0 )   b e g i n   a l u _ o u t _ T r a n s m i s s i o n   < =   0 ;   e n d  
                                 e l s e   b e g i n   a l u _ o u t _ T r a n s m i s s i o n   < =   1 ;   e n d  
               C M P _ P r e s s u r e :     i f ( d a t a _ 2 < = 9 ' h 0 f 0 )   b e g i n   a l u _ o u t _ P r e s s u r e   < =   0 ;   e n d  
                                 e l s e   b e g i n   a l u _ o u t _ P r e s s u r e   < =   1 ;   e n d  
             C M P _ O I L :     i f ( d a t a _ 2 < = 9 ' h 0 f 0 )   b e g i n   a l u _ o u t _ O I L   < =   0 ;   e n d  
                                 e l s e   b e g i n   a l u _ o u t _ O I L   < =   1 ;   e n d  
             C M P _ T e m p e r a t u r e :     i f ( d a t a _ 2 < = 9 ' h 0 f 0 )   b e g i n   a l u _ o u t _ t e m p e r a t u r e   < =   0 ;   e n d  
                                 e l s e   b e g i n   a l u _ o u t _ t e m p e r a t u r e   < =   1 ;   e n d  
             C M P _ b a t t e r y :     i f ( d a t a _ 2 < = 9 ' h 0 f 0 )   b e g i n   a l u _ o u t _ b a t t e r y   < =   0 ;   e n d  
                                 e l s e   b e g i n   a l u _ o u t _ b a t t e r y   < =   1 ;   e n d  
             d e f a u l t :   a l u _ o u t   =   0 ;  
         e n d c a s e  
 e n d m o d u l e  
  
  
 m o d u l e   C o n t r o l _ U n i t   (  
     L o a d _ R 0 ,   L o a d _ R 1 ,    
     L o a d _ R 2 ,   L o a d _ R 3 ,    
     L o a d _ P C ,   I n c _ P C ,    
     S e l _ B u s _ 1 _ M u x ,   S e l _ B u s _ 2 _ M u x ,  
     L o a d _ I R ,   L o a d _ A d d _ R ,   L o a d _ R e g _ Y ,   L o a d _ R e g _ Z ,    
     w r i t e ,   i n s t r u c t i o n ,   z e r o ,   c l k ,   r s t ) ;  
    
     p a r a m e t e r   w o r d _ s i z e   =   9 ,   o p _ s i z e   =   4 ,   s t a t e _ s i z e   =   4 ;  
     p a r a m e t e r   s r c _ s i z e   =   2 ,   d e s t _ s i z e   =   2 ,   S e l 1 _ s i z e   =   3 ,   S e l 2 _ s i z e   =   2 ;  
     / /   S t a t e   C o d e s  
     p a r a m e t e r   S _ i d l e   =   0 ,   S _ f e t 1   =   1 ,   S _ f e t 2   =   2 ,   S _ d e c   =   3 ;  
     p a r a m e t e r     S _ e x 1   =   4 ,   S _ r d 1   =   5 ,   S _ r d 2   =   6 ;      
     p a r a m e t e r   S _ w r 1   =   7 ,   S _ w r 2   =   8 ,   S _ b r 1   =   9 ,   S _ b r 2   =   1 0 ,   S _ h a l t   =   1 1 ;      
     / /   O p c o d e s  
     p a r a m e t e r   N O P   =   0 ,   A D D   =   1 ,   S U B   =   2 ,   A N D   =   3 ,   N O T   =   4 ;  
     p a r a m e t e r   R D     =   5 ,   W R   =     6 ,     B R   =     7 ,   B R Z   =   8 ;      
         p a r a m e t e r   C M P G a s   =   4 ' b 1 0 0 1 ;  
     p a r a m e t e r   C M P O i l   =   4 ' b 1 0 1 0 ;  
     p a r a m e t e r   C M P P r e s s u r e   =   4 ' b 1 0 1 1 ;  
     p a r a m e t e r   C M P T r a n s m i t t i o n   =   4 ' b 1 1 0 0 ;  
     p a r a m e t e r   C M P T e m p e r a t u r e   =   4 ' b 1 1 0 1 ;  
     p a r a m e t e r   C M P B a t t e r y   =   4 ' b 1 1 1 0 ;  
     / /   S o u r c e   a n d   D e s t i n a t i o n   C o d e s      
     p a r a m e t e r   R 0   =   0 ,   R 1   =   1 ,   R 2   =   2 ,   R 3   =   3 ;      
  
     o u t p u t   L o a d _ R 0 ,   L o a d _ R 1 ,   L o a d _ R 2 ,   L o a d _ R 3 ;  
     o u t p u t   L o a d _ P C ,   I n c _ P C ;  
     o u t p u t   [ S e l 1 _ s i z e - 1 : 0 ]   S e l _ B u s _ 1 _ M u x ;  
     o u t p u t   L o a d _ I R ,   L o a d _ A d d _ R ;  
     o u t p u t   L o a d _ R e g _ Y ,   L o a d _ R e g _ Z ;  
     o u t p u t   [ S e l 2 _ s i z e - 1 :   0 ]   S e l _ B u s _ 2 _ M u x ;  
     o u t p u t   w r i t e ;  
     i n p u t   [ w o r d _ s i z e - 1 :   0 ]   i n s t r u c t i o n ;  
     i n p u t   z e r o ;  
     i n p u t   c l k ,   r s t ;  
    
     r e g   [ s t a t e _ s i z e - 1 :   0 ]   s t a t e ,   n e x t _ s t a t e ;  
     r e g   L o a d _ R 0 ,   L o a d _ R 1 ,   L o a d _ R 2 ,   L o a d _ R 3 ,   L o a d _ P C ,   I n c _ P C ;  
     r e g   L o a d _ I R ,   L o a d _ A d d _ R ,   L o a d _ R e g _ Y ;  
     r e g   S e l _ A L U ,   S e l _ B u s _ 1 ,   S e l _ M e m ;  
     r e g   S e l _ R 0 ,   S e l _ R 1 ,   S e l _ R 2 ,   S e l _ R 3 ,   S e l _ P C ;  
     r e g   L o a d _ R e g _ Z ,   w r i t e ;  
     r e g   e r r _ f l a g ;  
  
     w i r e   [ o p _ s i z e - 1 : 0 ]   o p c o d e   =   i n s t r u c t i o n   [ w o r d _ s i z e - 1 :   w o r d _ s i z e   -   o p _ s i z e ] ;  
     w i r e   [ s r c _ s i z e - 1 :   0 ]   s r c   =   i n s t r u c t i o n   [ s r c _ s i z e   +   d e s t _ s i z e   - 1 :   d e s t _ s i z e ] ;  
     w i r e   [ d e s t _ s i z e - 1 : 0 ]   d e s t   =   i n s t r u c t i o n   [ d e s t _ s i z e   - 1 : 0 ] ;  
    
     / /   M u x   s e l e c t o r s  
     a s s i g n     S e l _ B u s _ 1 _ M u x [ S e l 1 _ s i z e - 1 : 0 ]   =   S e l _ R 0   ?   0 :  
 	 	 	 	   S e l _ R 1   ?   1 :  
 	 	 	 	   S e l _ R 2   ?   2 :  
 	 	 	 	   S e l _ R 3   ?   3 :  
 	 	 	 	   S e l _ P C   ?   4 :   3 ' b x ;     / /   3 - b i t s ,   s i z e d   n u m b e r  
  
     a s s i g n     S e l _ B u s _ 2 _ M u x [ S e l 2 _ s i z e - 1 : 0 ]   =   S e l _ A L U   ?   0 :  
 	 	 	 	   S e l _ B u s _ 1   ?   1 :  
 	 	 	 	   S e l _ M e m   ?   2 :   2 ' b x ;  
  
     a l w a y s   @   ( p o s e d g e   c l k   o r   n e g e d g e   r s t )   b e g i n :   S t a t e _ t r a n s i t i o n s  
         i f   ( r s t   = =   0 )   s t a t e   < =   S _ i d l e ;   e l s e   s t a t e   < =   n e x t _ s t a t e ;   e n d  
  
 / *     a l w a y s   @   ( s t a t e   o r   i n s t r u c t i o n   o r   z e r o )   b e g i n :     O u t p u t _ a n d _ n e x t _ s t a t e 	  
  
 N o t e :   T h e   a b o v e   e v e n t   c o n t r o l   e x p r e s s i o n   l e a d s   t o   i n c o r r e c t   o p e r a t i o n .     T h e   s t a t e   t r a n s i t i o n   c a u s e s   t h e   a c t i v i t y   t o   b e   e v a l u a t e d   o n c e ,   t h e n   t h e   r e s u l t i n g   i n s t r u c t i o n   c h a n g e   c a u s e s   i t   t o   b e   e v a l u a t e d   a g a i n ,   b u t   w i t h   t h e   r e s i d u a l   v a l u e   o f   o p c o d e .     O n   t h e   s e c o n d   p a s s   t h e   v a l u e   s e e n   i s   t h e   v a l u e   o p c o d e   h a d   b e f o r e   t h e   s t a t e   c h a n g e ,   w h i c h   r e s u l t s   i n   S e l _ P C   =   0   i n   s t a t e   3 ,   w h i c h   w i l l   c a u s e   a   r e t u r n   t o   s t a t e   1   a t   t h e   n e x t   c l o c k .     F i n a l l y ,   o p c o d e   i s   c h a n g e d ,   b u t   t h i s   d o e s   n o t   t r i g g e r   a   r e - e v a l u a t i o n   b e c a u s e   i t   i s   n o t   i n   t h e   e v e n t   c o n t r o l   e x p r e s s i o n .     S o ,   t h e   c a u t i o n   i s   t o   b e   s u r e   t o   u s e   o p c o d e   i n   t h e   e v e n t   c o n t r o l   e x p r e s s i o n .   T h a t   w a y ,   t h e   f i n a l   e x e c u t i o n   o f   t h e   b e h a v i o r   u s e s   t h e   v a l u e   o f   o p c o d e   t h a t   r e s u l t s   f r o m   t h e   s t a t e   c h a n g e ,   a n d   l e a d s   t o   t h e   c o r r e c t   v a l u e   o f   S e l _ P C .  
 * /    
  
     a l w a y s   @   ( s t a t e   o r   o p c o d e   o r   z e r o )   b e g i n :   O u t p u t _ a n d _ n e x t _ s t a t e    
         S e l _ R 0   =   0 ;   	 S e l _ R 1   =   0 ;           	 S e l _ R 2   =   0 ;         	 S e l _ R 3   =   0 ;           	 S e l _ P C   =   0 ;  
         L o a d _ R 0   =   0 ;   	 L o a d _ R 1   =   0 ;   	 L o a d _ R 2   =   0 ;   	 L o a d _ R 3   =   0 ; 	 L o a d _ P C   =   0 ;  
  
         L o a d _ I R   =   0 ; 	 L o a d _ A d d _ R   =   0 ; 	 L o a d _ R e g _ Y   =   0 ; 	 L o a d _ R e g _ Z   =   0 ;  
         I n c _ P C   =   0 ;    
         S e l _ B u s _ 1   =   0 ;    
         S e l _ A L U   =   0 ;    
         S e l _ M e m   =   0 ;    
         w r i t e   =   0 ;    
         e r r _ f l a g   =   0 ; 	 / /   U s e d   f o r   d e - b u g   i n   s i m u l a t i o n 	 	  
          
         n e x t _ s t a t e   =   s t a t e ;  
          
  
           c a s e     ( s t a t e ) 	 S _ i d l e : 	 	 n e x t _ s t a t e   =   S _ f e t 1 ;              
 S _ f e t 1 : 	 	 b e g i n               	     	     	  
     n e x t _ s t a t e   =   S _ f e t 2 ;    
             	     	     	 	     S e l _ P C   =   1 ;  
             	     	     	 	     S e l _ B u s _ 1   =   1 ;  
             	     	       	 	     L o a d _ A d d _ R   =   1 ;    
         	 	 	 	 e n d  
             	 	 S _ f e t 2 : 	 	 b e g i n   	 	  
     n e x t _ s t a t e   =   S _ d e c ;    
     S e l _ M e m   =   1 ;  
             	     	     	 	     L o a d _ I R   =   1 ;    
             	     	     	 	     I n c _ P C   =   1 ;  
         	 	 	 	 e n d  
  
             	 	 S _ d e c :     	   	 c a s e     ( o p c o d e )    
             	 	   	 	     N O P :   n e x t _ s t a t e   =   S _ f e t 1 ;  
 	 	     	 	     A D D ,   S U B ,   A N D :   b e g i n  
   	 	         	 	         n e x t _ s t a t e   =   S _ e x 1 ;  
 	 	         	 	         S e l _ B u s _ 1   =   1 ;  
 	 	         	 	         L o a d _ R e g _ Y   =   1 ;  
 	 	           	 	         c a s e     ( s r c )  
 	 	             	 	             R 0 :   	 	 S e l _ R 0   =   1 ;    
 	 	             	 	             R 1 :   	 	 S e l _ R 1   =   1 ;    
 	 	             	 	             R 2 :   	 	 S e l _ R 2   =   1 ;  
 	 	             	 	             R 3 :   	 	 S e l _ R 3   =   1 ;    
 	 	             	 	             d e f a u l t   :   	 e r r _ f l a g   =   1 ;  
 	 	         	 	         e n d c a s e        
     e n d   / /   A D D ,   S U B ,   A N D  
  
 	 	 	   	     N O T , C M P G a s ,   C M P O i l , C M P P r e s s u r e ,   C M P T r a n s m i t t i o n , C M P T e m p e r a t u r e , C M P B a t t e r y :   b e g i n  
 	 	 	         	         n e x t _ s t a t e   =   S _ f e t 1 ;  
 	 	 	         	         L o a d _ R e g _ Z   =   1 ;  
 	 	 	         	         S e l _ B u s _ 1   =   1 ;    
 	 	 	         	         S e l _ A L U   =   1 ;    
 	 	   	           	         c a s e     ( s r c )  
 	 	 	             	             R 0 :   	 	 S e l _ R 0   =   1 ; 	 	 	              
             	 	 	 	             R 1 :   	 	 S e l _ R 1   =   1 ;  
 	 	 	             	             R 2 :   	 	 S e l _ R 2   =   1 ; 	 	 	              
   	 	 	             	             R 3 :   	 	 S e l _ R 3   =   1 ;    
 	 	 	             	             d e f a u l t   :   	 e r r _ f l a g   =   1 ;  
 	 	 	         	         e n d c a s e        
     	 	 	           	         c a s e     ( d e s t )  
 	 	 	             	             R 0 :   	 	 L o a d _ R 0   =   1 ;    
 	 	 	             	             R 1 :   	 	 L o a d _ R 1   =   1 ; 	 	 	              
             	 	 	 	             R 2 :   	 	 L o a d _ R 2   =   1 ;  
 	 	 	             	             R 3 :   	 	 L o a d _ R 3   =   1 ; 	 	 	              
             	 	 	 	             d e f a u l t :   	 e r r _ f l a g   =   1 ;  
 	 	 	         	         e n d c a s e        
     e n d   / /   N O T  
     	 	 	 	      
     R D :   b e g i n  
 	 	 	         	         n e x t _ s t a t e   =   S _ r d 1 ;  
 	 	 	         	         S e l _ P C   =   1 ;   S e l _ B u s _ 1   =   1 ;   L o a d _ A d d _ R   =   1 ;    
     e n d   / /   R D  
  
 	 	 	     	     W R :   b e g i n  
 	 	 	         	         n e x t _ s t a t e   =   S _ w r 1 ;  
 	 	 	         	         S e l _ P C   =   1 ;   S e l _ B u s _ 1   =   1 ;   L o a d _ A d d _ R   =   1 ;    
     e n d     / /   W R  
  
 	 	 	     	     B R :   b e g i n    
 	 	 	         	         n e x t _ s t a t e   =   S _ b r 1 ;      
         S e l _ P C   =   1 ;   S e l _ B u s _ 1   =   1 ;   L o a d _ A d d _ R   =   1 ;    
 	 	 	         	     e n d     / /   B R  
 	  
     	 	 	 	     B R Z :   i f   ( z e r o   = =   1 )   b e g i n  
 	 	 	         	         n e x t _ s t a t e   =   S _ b r 1 ;    
         S e l _ P C   =   1 ;   S e l _ B u s _ 1   =   1 ;   L o a d _ A d d _ R   =   1 ;    
 	 	 	         	     e n d   / /   B R Z  
 	 	 	     	     e l s e   b e g i n    
         n e x t _ s t a t e   =   S _ f e t 1 ;    
         I n c _ P C   =   1 ;    
     e n d  
      
    
                 	 	     	 	     d e f a u l t   :   n e x t _ s t a t e   =   S _ h a l t ;  
 	 	 	 	 e n d c a s e     / /   ( o p c o d e )  
  
         	             	 S _ e x 1 : 	 	 b e g i n    
     	 	 	     	     n e x t _ s t a t e   =   S _ f e t 1 ;  
 	 	 	     	     L o a d _ R e g _ Z   =   1 ;  
 	 	 	     	     S e l _ A L U   =   1 ;    
 	 	   	       	     c a s e     ( d e s t )  
     	         	 	         	         R 0 :   b e g i n   S e l _ R 0   =   1 ;   L o a d _ R 0   =   1 ;   e n d  
 	 	 	         	         R 1 :   b e g i n   S e l _ R 1   =   1 ;   L o a d _ R 1   =   1 ;   e n d  
 	 	 	         	         R 2 :   b e g i n   S e l _ R 2   =   1 ;   L o a d _ R 2   =   1 ;   e n d  
 	 	 	         	         R 3 :   b e g i n   S e l _ R 3   =   1 ;   L o a d _ R 3   =   1 ;   e n d  
 	 	 	         	         d e f a u l t   :   e r r _ f l a g   =   1 ;    
 	 	 	       	     e n d c a s e      
 	 	 	 	 e n d    
  
         	             	 S _ r d 1 : 	 	 b e g i n    
     n e x t _ s t a t e   =   S _ r d 2 ;  
 	 	 	     	     S e l _ M e m   =   1 ;  
 	 	 	     	     L o a d _ A d d _ R   =   1 ;    
 	 	 	     	     I n c _ P C   =   1 ;  
 	 	 	 	 e n d  
  
         	             	 S _ w r 1 :   	 	 b e g i n  
 	 	 	     	     n e x t _ s t a t e   =   S _ w r 2 ;  
 	 	 	     	     S e l _ M e m   =   1 ;  
 	 	 	     	     L o a d _ A d d _ R   =   1 ;    
 	 	 	     	     I n c _ P C   =   1 ;  
 	 	 	 	 e n d    
  
             	 	 S _ r d 2 : 	 	 b e g i n    
     	 	 	     	     n e x t _ s t a t e   =   S _ f e t 1 ;  
 	 	 	     	     S e l _ M e m   =   1 ;  
 	 	   	       	     c a s e     ( d e s t )    
         	 	 	         	         R 0 :   	 	 L o a d _ R 0   =   1 ;    
 	 	   	         	         R 1 :   	 	 L o a d _ R 1   =   1 ;    
 	 	   	         	         R 2 :   	 	 L o a d _ R 2   =   1 ;    
 	 	   	         	         R 3 :   	 	 L o a d _ R 3   =   1 ;    
 	 	 	         	         d e f a u l t   :   	 e r r _ f l a g   =   1 ;  
 	 	 	     	     e n d c a s e      
 	 	 	 	 e n d  
  
         	             	 S _ w r 2 : 	 	 b e g i n    
           	 	 	     	     n e x t _ s t a t e   =   S _ f e t 1 ;  
 	 	 	     	     w r i t e   =   1 ;  
 	 	   	     	     c a s e     ( s r c )  
         	 	 	         	         R 0 :   	 	 S e l _ R 0   =   1 ; 	 	   	          
         	 	 	 	         R 1 :   	 	 S e l _ R 1   =   1 ; 	 	   	          
       	 	 	 	         R 2 :   	 	 S e l _ R 2   =   1 ;   	 	   	          
       	 	 	 	         R 3 :   	 	 S e l _ R 3   =   1 ; 	 	 	          
         	 	 	 	         d e f a u l t   :   	 e r r _ f l a g   =   1 ;  
 	 	 	     	     e n d c a s e      
 	 	 	 	 e n d  
  
         	             	 S _ b r 1 : 	 	 b e g i n   n e x t _ s t a t e   =   S _ b r 2 ;   S e l _ M e m   =   1 ;   L o a d _ A d d _ R   =   1 ;   e n d  
         	             	 S _ b r 2 : 	 	 b e g i n   n e x t _ s t a t e   =   S _ f e t 1 ;   S e l _ M e m   =   1 ;   L o a d _ P C   =   1 ;   e n d  
         	             	 S _ h a l t :     	 	 n e x t _ s t a t e   =   S _ h a l t ;  
         	             	  
 	 	 d e f a u l t : 	 	 n e x t _ s t a t e   =   S _ i d l e ;  
           e n d c a s e          
     e n d  
 e n d m o d u l e  
  
  
 m o d u l e   M e m o r y _ U n i t   ( d a t a _ o u t ,   d a t a _ i n ,   a d d r e s s ,   c l k ,   w r i t e ) ;  
     p a r a m e t e r   w o r d _ s i z e   =   9 ;  
     p a r a m e t e r   m e m o r y _ s i z e   =   5 1 2 ;  
  
     o u t p u t   [ w o r d _ s i z e - 1 :   0 ]   d a t a _ o u t ;  
     i n p u t   [ w o r d _ s i z e - 1 :   0 ]   d a t a _ i n ;  
     i n p u t   [ w o r d _ s i z e - 1 :   0 ]   a d d r e s s ;  
     i n p u t   c l k ,   w r i t e ;  
     r e g   [ w o r d _ s i z e - 1 :   0 ]   m e m o r y   [ m e m o r y _ s i z e - 1 :   0 ] ;  
  
     a s s i g n   d a t a _ o u t   =   m e m o r y [ a d d r e s s ] ;  
  
     a l w a y s   @   ( p o s e d g e   c l k )  
         i f   ( w r i t e )   m e m o r y [ a d d r e s s ]   =   d a t a _ i n ;  
 e n d m o d u l e  
  
 